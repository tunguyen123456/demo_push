library verilog;
use verilog.vl_types.all;
entity Lab_06_vlg_vec_tst is
end Lab_06_vlg_vec_tst;
