library verilog;
use verilog.vl_types.all;
entity up_down_vlg_check_tst is
    port(
        Y0              : in     vl_logic;
        Y1              : in     vl_logic;
        Y2              : in     vl_logic;
        Y3              : in     vl_logic;
        Y4              : in     vl_logic;
        Y5              : in     vl_logic;
        Y6              : in     vl_logic;
        Y7              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end up_down_vlg_check_tst;
