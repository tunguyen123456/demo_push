library verilog;
use verilog.vl_types.all;
entity up_down is
    port(
        Y3              : out    vl_logic;
        D               : in     vl_logic;
        E               : in     vl_logic;
        LOAD            : in     vl_logic;
        I3              : in     vl_logic;
        I2              : in     vl_logic;
        I1              : in     vl_logic;
        I0              : in     vl_logic;
        CLK             : in     vl_logic;
        Y2              : out    vl_logic;
        Y7              : out    vl_logic;
        I7              : in     vl_logic;
        I6              : in     vl_logic;
        I5              : in     vl_logic;
        I4              : in     vl_logic;
        Y6              : out    vl_logic;
        Y0              : out    vl_logic;
        Y1              : out    vl_logic;
        Y4              : out    vl_logic;
        Y5              : out    vl_logic
    );
end up_down;
