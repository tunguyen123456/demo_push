library verilog;
use verilog.vl_types.all;
entity Lab_06_KhongCuBo_vlg_check_tst is
    port(
        O               : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end Lab_06_KhongCuBo_vlg_check_tst;
